��   A��A��*SYST�EM*��V9.3�0259 9/�14/2023 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1 N � �CLo: �� �AX{  �$PS_�TI����TIME ��J� _CMD,��"FB�VS �&�CL_OV�� F�RMZ�$DED�X�$NA� %��CURL�W����TCK5�wFMSV�M_LIF	��`;8G:w$�A9_0M:_��=�93x6W� |�"�PCCOM���FB� M�0�M7AL_�ECIr�PL!�"DTYk�R_�"�5L#�1EN�DD��o1� �5M� b��PL� W � � $STAL#TRGQ_M��0KN}FS� �HY�J� |G�I�JI�JI�E#3�AnCuB�A���$��ASS> ����	Q�����@V�ERSI� W�  1���$S 1'X� ���N ���n_Y_�_}U���8��)�
�i]��_��X_ �_�_�_x_�Q.g;o�S�QTico�Q��� �ᩁ�Fm�i}�do_�o�f`o��o�o�o�o!�dw@
Mv @
8 �o�k���d�� ��� �2�D�V�h� z�������ԏ��� 
��.�@��{	Ue�s�8]���T  2�ğ ֟�����0�B�T�f��R��������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬϾ�������� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n������<���������&��8�J�\�n������|( ����������2 /hS�w�� ���
�.R =v�o���� ��/*//N/9/r/ +�/�/�/�/�/�/W/  ?&??J?5?n?�}�� �?�?�?�?�?�?OO /OAOSOeOwO�O���O �O�O�O�O_R��Ov� (_^_���_�_�_�_�_ �_�_oo'or�Ko]o oo�o�o�o�o�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _���Ho������˯ݯ ���%�7�I�[�{� nPLQ����`?����տ �������/��S�>��w�bϛφϘ��� ��$FMS_GRP� 1mU� ���T���O�r�Pr?7�Qu�h�ϻ��?�&AE���B��=]�0<߻�6!}V�A��ω�t߭ߘ�A�  ���ߠ����+���O�:�s���Ymn�Z�|qn���}� ���j����f����+�=�x�% � ot a programH�z��� "������������P� b�3����iT�x ����A�$ �H3l~��� i��/�2/D/ �h/z/��//�/�/ �/�/K/?.?�/�/d? �/�?s?�?�??�?�? G?�?*OONO9OrO�O �?�O�OO�OYO__ �O8_�O\_n_�O#_�_ _�_�_�_�_Q_"o4o �_�_joUo�oyo�o�o o�o�oMo�oBT ?x�o��c� _��,�>��b�t� �)�����Ώ���� W�(�:���^�ُ���� ����ܟ�A���$� ��H�3�l�~�џ���� �i��կ���2�D� ��h�z�ͯ���¿Կ ����K��.ρ��d� ߿��sϬϾ������ Gϩ�*��N�9�r߄�p�Ϩߺ�e����� ��e����*��N�9� r��o�������� ����&��J�5�n��8_��� �����V�������-��23�456789010QY~�����ц ��������� ����R�vd ����8�/ /</*/`/r/��/� �x/J/�/?�/&?|/ �/_?�/�/�??�?�? �?�?B?O%Ox?�?XO FO|OjO�O�OO�O,O >O�O�O_B_0_f_�O �O�_�O_�_P_�_�_ o,o�_Soeo�_o�o �o�o�o�o�oHolo ~o�o�oL�p��o �2D��6�$� F�l�������Z�؏ Ə��� �2���Y��� ��8�
������<� N��r���R�Пv�d� �����ӯ�8���� �<�*�`�r�ȯ��� ��x�J�̿��&�|� ��_ϲ�Ŀ��϶Ϥ� ����B��%�x���X� F�|�jߠ߲����,� >߸ߊ��B�0�f�x뀇��ߟ���������$PLCL_GR�P 1]��� p?�  �"���E�i� T���x����������� ��/ �bL� ,������ +O:s^�� x�p